netcdf tpoce_MED-12_ERA5_evaluation_r1i1p1f1_CNRM-MF_CNRM-RCSM6B-SN_v1-r1_mon_198803-198803 {
dimensions:
	axis_nbounds = 2 ;
	x = 567 ;
	y = 264 ;
	deptht = 75 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float nav_lat(y, x) ;
		nav_lat:standard_name = "latitude" ;
		nav_lat:long_name = "Latitude" ;
		nav_lat:units = "degrees_north" ;
	float nav_lon(y, x) ;
		nav_lon:standard_name = "longitude" ;
		nav_lon:long_name = "Longitude" ;
		nav_lon:units = "degrees_east" ;
	float deptht(deptht) ;
		deptht:name = "deptht" ;
		deptht:long_name = "Vertical T levels" ;
		deptht:units = "m" ;
		deptht:positive = "down" ;
		deptht:bounds = "deptht_bounds" ;
	float deptht_bounds(deptht, axis_nbounds) ;
		deptht_bounds:units = "m" ;
	double time(time) ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:long_name = "Time axis" ;
		time:calendar = "gregorian" ;
		time:units = "days since 1900-01-01 00:00:00" ;
		time:time_origin = "1900-01-01 00:00:00" ;
		time:bounds = "time_bounds" ;
	double time_bounds(time, axis_nbounds) ;
	float tpoce(time, deptht, y, x) ;
		tpoce:standard_name = "sea_water_potential_temperature" ;
		tpoce:long_name = "Sea Water Potential Temperature" ;
		tpoce:units = "degC" ;
		tpoce:online_operation = "average" ;
		tpoce:cell_methods = "time: mean" ;
		tpoce:interval_operation = "720 s" ;
		tpoce:interval_write = "1 month" ;
		tpoce:_FillValue = 1.e+20f ;
		tpoce:missing_value = 1.e+20f ;
		tpoce:coordinates = "nav_lat nav_lon" ;
		tpoce:description = "None" ;
		tpoce:history = "none" ;
		tpoce:cell_measures = "area: areacello" ;

// global attributes:
		:name = "/scratch/work/sevault/CNRM-RCSM6B/RCSM6B-ERA5.2/outputs/19880101/tpoce_MED-12_ERA5_evaluation_r1i1p1f1_CNRM-MF_CNRM-RCSM6B-SN_v1-r1_mon_%start_date%-%end_date%" ;
		:description = "Created by xios" ;
		:creation_date = "2024-03-29T07:43:23Z" ;
		:tracking_id = "hdl:21.14103/227c3a13-dde3-4b47-987e-3d7e0120cae1" ;
		:title = "CNRM-RCSM6B-SN model output prepared for CORDEX-CMIP6 / evaluation simulation driven by ERA5, evaluation, r1i1p1f1" ;
		:Conventions = "CF-1.10" ;
		:activity_id = "RCM" ;
		:comment = "CORDEX MED-12 CNRM-RCSM6B-SN L91." ;
		:contact = "contact.aladin-cordex@meteo.fr" ;
		:dr2xml_version = "3.0" ;
		:domain = "MED-12" ;
		:domain_id = "MED-12" ;
		:driving_experiment = "ERA5, evaluation, r1i1p1f1" ;
		:driving_experiment_id = "evaluation" ;
		:driving_institution_id = "ECMWF" ;
		:driving_source_id = "ERA5" ;
		:driving_variant_label = "r1i1p1f1" ;
		:experiment_id = "evaluation" ;
		:external_variables = "areacello" ;
		:frequency = "mon" ;
		:further_info_url = "http://www.umr-cnrm.fr/" ;
		:history = "none" ;
		:institution = "CNRM (Centre National de Recherches Meteorologiques) - Météo France, Toulouse, France" ;
		:institution_id = "CNRM-MF" ;
		:license = "CORDEX model data produced by CNRM-MF is licensed under a Creative Commons Attribution 4.0 International License (https://creativecommons.org/licenses). Consult (...) for terms of use governing CORDEX output, including citation requirements and proper acknowledgment. The data producers and data providers make no warranty, either express or implied, including, but not limited to, warranties of merchantability and fitness for a particular purpose. All liabilities arising from the supply of the information (including any liability arising in negligence) are excluded to the fullest extent permitted by law." ;
		:mip_era = "CMIP6" ;
		:native_resolution = "8 km" ;
		:product = "model-output" ;
		:project_id = "CORDEX" ;
		:realm = "ocean" ;
		:references = "Nabat, P., Somot, S., Cassou, C., Mallet, M., Michou, M., Bouniol, D., Decharme, B., Druge, T., Roehrig, R. and Saint-Martin, D. (2020): Modulation of radiative aerosols effects by atmospheric circulation over the Euro-Mediterranean region, Atmos. Chem. Phys., 20, 8315-8349, doi:10.5194/acp-20-8315-2020." ;
		:source = "CNRM-ALADIN64E1" ;
		:source_id = "CNRM-ALADIN64E1" ;
		:source_type = "AORCM AER" ;
		:variable_id = "tpoce" ;
		:version_realisation = "v1-r1" ;
		:CMIP6_CV_version = "cv=6.2.3.0-7-g2019642" ;
		:EXPID = "RCSM6B-ERA5.2" ;
		:dr2xml_md5sum = "fdee7e9a1c0c1c2cb709a65fb5c920d5" ;
		:xios_commit = "1442-shuffle" ;
}
